/******************************************************************************
 * (C) Copyright 2014 AMIQ Consulting
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * NAME:        amiq_hello_world_import_functions.svh
 * PROJECT:     amiq_hello_world
 * Description: Forward declaration for all functions imported from DPI-C
 *******************************************************************************/
 
`ifndef __amiq_hello_world_import_functions
    `define __amiq_hello_world_import_functions

// Initialize the octave API
import "DPI-C" function void initialize_octave();

// Hello world example C function
import "DPI-C" function void c_hello_world();

`endif
